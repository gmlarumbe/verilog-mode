module align_param # (
parameter PARAM_1 = 0,
parameter PARAMETER_2 = 1
);

localparam LOCAL_1 = 1;
localparam LOCAL_LONG = 2;
localparam LOCAL_MULTILINE = 3,
LOCAL2 = 4,
LOCAL_LONG3 = 5;

endmodule


// Local Variables:
// verilog-align-param-expr: nil
// End:
