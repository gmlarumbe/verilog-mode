interface class ic;
   // ...
endclass
   // this should indent to left margin, but indents one stop to right
