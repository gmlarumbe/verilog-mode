module foo (input logic [7:0] in1,
            input logic       in2,
            custom_type       type1,
            output logic      out,
            custom_type       type2
            );
   
   logic [7:0] signal1;
   logic       signal2;
   custom_type type3;
   
endmodule

// Local Variables:
// eval: (setq verilog-declaration-typedef-words '("custom_type"))
// End:
